// Hello World in Verilog
module hello_world;

  initial begin
    // Display "Hello, World!" to the console
    $display("Hello, World!");
    // End the simulation
    $finish;
  end

endmodule
